library verilog;
use verilog.vl_types.all;
entity SSD1306_VHDLImplementation_vlg_vec_tst is
end SSD1306_VHDLImplementation_vlg_vec_tst;
