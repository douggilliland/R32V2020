-- Timer/Counter Unit
-- Contains three counters
--		System clock counter (when 50 MHz clock, counts are in 20 nS increments)
--		microsecond counter (accuracy is +/- 1 uS)
--		millisecond counter (accuracy is +/- 1 mSec)
--		Elapsed time counter (accuracy is +/- 1 CPU clock)

library ieee;
use ieee.std_logic_1164.all;
use  IEEE.STD_LOGIC_ARITH.all;
use  IEEE.STD_LOGIC_UNSIGNED.all;
library work;
use work.R32V2020_Pkg.all;

entity Timer_Unit is
	port(
		n_reset						: in std_logic := '1';
		i_CLOCK_50					: in std_logic := '1';
		i_OneHotState				: in std_logic_vector(3 downto 0) := "0000";
		-- Peripheral Memory Mapped Space Address/Data/Control lines
 		i_peripheralWrStrobe		: in std_logic := '1';
		i_peripheralAddress		: in std_logic_vector(31 downto 0) := x"00000000";
		i_dataToTimers				: in std_logic_vector(31 downto 0) := x"00000000";
		o_dataFromTimers			: out std_logic_vector(31 downto 0) := x"00000000"
		);
	end Timer_Unit;

	architecture struct of Timer_Unit is

	--attribute syn_keep: boolean;
	-- Peripheral Signals
	signal w_ElapsedTimeCount		:	std_logic_vector(31 downto 0);
	signal q_MicrosecondScaler		: 	std_logic_vector(5 downto 0);
	signal q_MicrosecondCounter	: 	std_logic_vector(31 downto 0);
	signal q_MillisecondScaler		: 	std_logic_vector(10 downto 0);
	signal q_MillisecondCounter	: 	std_logic_vector(31 downto 0);
	signal q_CPUCycleCounter		: 	std_logic_vector(31 downto 0);

begin
	o_dataFromTimers <= 
	w_ElapsedTimeCount 	when i_peripheralAddress(2 downto 0) = "000" else	-- Counts in FPGA clock ticks (50 MHz for most FPGAs)
	q_MicrosecondCounter when i_peripheralAddress(2 downto 0) = "001" else	-- Counts in uSecs
	q_MillisecondCounter when i_peripheralAddress(2 downto 0) = "010" else	-- Counts in mSecs
	q_CPUCycleCounter 	when i_peripheralAddress(2 downto 0) = "011" else	-- Counts CPU instructions
	x"00000000";

	-- Elapsed Time Counter
	ETC : entity work.COUNT_32
	Port map (
		clk 		=> i_CLOCK_50,
		clr 		=> not n_reset,
		d   		=> x"00000000",
		enable	=> '1',
		inc 		=> '1',
		dec		=> '0',
		q   		=> w_ElapsedTimeCount
	);
	
	process (i_CLOCK_50, n_reset)
	begin
		if (n_reset='0') then
			q_MicrosecondScaler 		<= (others => '0');
			q_MicrosecondCounter 	<= (others => '0');
			q_MillisecondScaler		<= (others => '0');
			q_MillisecondCounter 	<= (others => '0');
			q_CPUCycleCounter			<= (others => '0');
		elsif(rising_edge(i_CLOCK_50)) then
			if (i_OneHotState(0) = '1') then 
				q_CPUCycleCounter <= q_CPUCycleCounter + 1;
			end if;
			if (q_MicrosecondScaler < 49) then
				q_MicrosecondScaler <= q_MicrosecondScaler + 1;
			else	-- Microsecond terminal count
				q_MicrosecondScaler <= (others => '0');
				q_MicrosecondCounter <= q_MicrosecondCounter + 1;
				if (q_MillisecondScaler < 999) then	-- millisecond scaler
					q_MillisecondScaler <= q_MillisecondScaler + 1;
				else
					q_MillisecondScaler <= (others => '0');
					q_MillisecondCounter <= q_MillisecondCounter + 1;
				end if;
			end if;
			
		end if;
	end process;
	
end struct;
